`include "light_package.sv"
`include "traffic_light_controller.sv"