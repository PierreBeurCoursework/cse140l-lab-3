`include "lab3_part2_tb_enum.sv"