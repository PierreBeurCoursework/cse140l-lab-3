`include "light_package.sv"
`include "traffic_light_controller_starter_RRH.sv"