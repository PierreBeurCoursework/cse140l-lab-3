`include "lab3_part1_tb_enum.sv"